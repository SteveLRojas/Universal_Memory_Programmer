`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   14:44:11 06/15/2022
// Design Name:   Nexys2_programmer
// Module Name:   /home/ise/VM_share/Nexys2_programmer/testbench.v
// Project Name:  Nexys2_programmer
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: Nexys2_programmer
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module testbench;

	// Inputs
	reg clk;
	reg [3:0] button;
	wire rxd;
	reg flash_sts;

	// Outputs
	wire [7:0] led;
	wire txd;
	wire [22:0] flash_a;
	wire flash_we_n;
	wire flash_reset_n;
	wire flash_ce_n;
	wire flash_oe_n;
	wire psram_ce_n;
	wire [3:0] seg_sel;
	wire [7:0] hex_out;

	// Bidirs
	wire ps2_data;
	wire ps2_clk;
	wire [15:0] flash_d;
	
	pullup(ps2_data);
	pullup(ps2_clk);
	pullup(flash_d[0]);
	pullup(flash_d[1]);
	pullup(flash_d[2]);
	pullup(flash_d[3]);
	pullup(flash_d[4]);
	pullup(flash_d[5]);
	pullup(flash_d[6]);
	pullup(flash_d[7]);
	
	//internal signals
	wire[15:0] hex_indicators;
	wire[15:0] led_indicators;
	
	wire[15:0] IO_address;
	wire[15:0] from_cpu;
	wire[15:0] IO_to_cpu;
	wire IO_wren;
	wire IO_ren;
	wire L_en;
	wire H_en;

	// Instantiate the Unit Under Test (UUT)
	Nexys2_programmer uut (
		.clk(clk), 
		.button(button),
		.switch(2'b10),
		.led(led), 
		.rxd(rxd), 
		.txd(txd), 
		.ps2_data(ps2_data), 
		.ps2_clk(ps2_clk), 
		.shared_a(flash_a), 
		.shared_d(flash_d),
		.shared_oe_n(flash_oe_n),
		.shared_we_n(flash_we_n), 
		.flash_ce_n(flash_ce_n),
		.flash_reset_n(flash_reset_n), 
		.flash_sts(flash_sts), 
		.psram_ce_n(psram_ce_n),
		.psram_adv_n(),
		.psram_cre(),
		.psram_clk(),
		.psram_lb_n(),
		.psram_ub_n(),
		.seg_sel(seg_sel), 
		.hex_out(hex_out)
	);
	
	assign hex_indicators = uut.hex_indicators;
	assign led_indicators = uut.led_indicators;
	
	assign IO_address = uut.IO_address;
	assign from_cpu = uut.from_cpu;
	assign IO_to_cpu = uut.IO_to_cpu;
	assign IO_wren = uut.IO_wren;
	assign IO_ren = uut.IO_ren;
	assign L_en = uut.L_en;
	assign H_en = uut.H_en;
	
	//test inputs from PC
	reg[7:0] test_inputs[0:31];
	reg[4:0] test_index;
	reg test_tx_req;
	wire test_tx_ready;
	wire test_rx_ready;
	reg test_tx_busy;
	wire[7:0] test_tx_data;
	wire[7:0] test_rx_data;

	assign test_tx_data = test_inputs[test_index];

	UART test_UART(
				.clk(clk),
				.reset(button[0]),
				.tx_req(test_tx_req),
				.tx_data(test_tx_data),
				.rx(txd),
				.tx(rxd),
				.rx_data(test_rx_data),
				.tx_ready(test_tx_ready),
				.rx_ready(test_rx_ready));

	always @(posedge clk)
	begin
		test_tx_req <= 1'b0;
		if(button[0])
		begin
			test_tx_busy <= 1'b0;
			test_index <= 5'h0;
		end
		else
		begin
			if(test_tx_req)
				test_tx_busy <= 1'b1;
			if(test_tx_ready)
				test_tx_busy <= 1'b0;
			if(~test_tx_busy & (test_index != 5'h1f))
				test_tx_req <= 1'b1;
			if(test_tx_ready & (test_index != 5'h1f))
				test_index <= test_index + 5'h01;
		end
	end
	
	always
	begin
		#10 clk = ~clk;
	end

	initial begin
		// Initialize Inputs
		test_inputs[0] = 8'hde;
		test_inputs[1] = 8'had;
		test_inputs[2] = 8'hbe;
		test_inputs[3] = 8'hef;
		
		test_inputs[4] = 8'h01;
		
		test_inputs[5] = 8'h00;
		test_inputs[6] = 8'h00;
		test_inputs[7] = 8'h00;
		test_inputs[8] = 8'h10;
		
		test_inputs[9] = 8'h64;
		test_inputs[10] = 8'h65;
		test_inputs[11] = 8'h72;
		test_inputs[12] = 8'h67;
		test_inputs[13] = 8'h20;
		test_inputs[14] = 8'h77;
		test_inputs[15] = 8'h61;
		test_inputs[16] = 8'h73;
		test_inputs[17] = 8'h20;
		test_inputs[18] = 8'h68;
		test_inputs[19] = 8'h65;
		test_inputs[20] = 8'h72;
		test_inputs[21] = 8'h65;
		test_inputs[22] = 8'h2e;
		test_inputs[23] = 8'hde;
		test_inputs[24] = 8'had;
		test_inputs[25] = 8'hbe;
		test_inputs[26] = 8'hef;
		test_inputs[27] = 8'hde;
		test_inputs[28] = 8'had;
		test_inputs[29] = 8'hbe;
		test_inputs[30] = 8'hef;
		test_inputs[31] = 8'hde;
		
		clk = 0;
		flash_sts = 1'b1;
		button = 4'h1;

		// Wait 100 ns for global reset to finish
		#200 button = 4'h0;
        
		// Add stimulus here

	end
      
endmodule

